library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity inst_rom16 is
  port (
    address : in  std_logic_vector(7 downto 0);
    q       : out std_logic_vector(15 downto 0)
  );
end entity;

architecture rtl of inst_rom16 is
  type rom_t is array (0 to 255) of std_logic_vector(15 downto 0);
  constant rom : rom_t := (
    0   => x"5204",
    1   => x"7210",
    2   => x"5307",
    3   => x"7320",
    4   => x"53FD",
    5   => x"7321",
    6   => x"530C",
    7   => x"7322",
    8   => x"5300",
    9   => x"7323",
    10  => x"5300",
    11  => x"5120",
    12  => x"6600",
    13  => x"0EC2",
    14  => x"5501",
    15  => x"6600",
    16  => x"0EC2",
    17  => x"5501",
    18  => x"6600",
    19  => x"0EC2",
    20  => x"5501",
    21  => x"6600",
    22  => x"0EC2",
    23  => x"7311",
    24  => x"5200",
    25  => x"7213",
    26  => x"6313",
    27  => x"5203",
    28  => x"8E16",
    29  => x"5203",
    30  => x"0B83",
    31  => x"7215",
    32  => x"5200",
    33  => x"7214",
    34  => x"5120",
    35  => x"6600",
    36  => x"6701",
    37  => x"AB01",
    38  => x"8002",
    39  => x"7700",
    40  => x"7601",
    41  => x"5501",
    42  => x"6214",
    43  => x"5A01",
    44  => x"7214",
    45  => x"6315",
    46  => x"9BF4",
    47  => x"6213",
    48  => x"5A01",
    49  => x"7213",
    50  => x"B01A",
    51  => x"5120",
    52  => x"5300",
    53  => x"6600",
    54  => x"0EC2",
    55  => x"5501",
    56  => x"6600",
    57  => x"0EC2",
    58  => x"5501",
    59  => x"6600",
    60  => x"0EC2",
    61  => x"5501",
    62  => x"6600",
    63  => x"0EC2",
    64  => x"7312",
    65  => x"6211",
    66  => x"6312",
    67  => x"8B01",
    68  => x"B061",
    69  => x"5120",
    70  => x"6600",
    71  => x"6701",
    72  => x"0EC7",
    73  => x"9C17",
    74  => x"5501",
    75  => x"6600",
    76  => x"6701",
    77  => x"0EC7",
    78  => x"9C12",
    79  => x"5501",
    80  => x"6600",
    81  => x"6701",
    82  => x"0EC7",
    83  => x"9C0D",
    84  => x"6212",
    85  => x"4B0F",
    86  => x"5101",
    87  => x"0DC4",
    88  => x"0985",
    89  => x"0EC0",
    90  => x"0DC6",
    91  => x"0DC3",
    92  => x"0EC1",
    93  => x"220A",
    94  => x"3AAA",
    95  => x"1800",
    96  => x"C000",
    97  => x"220E",
    98  => x"3AEE",
    99  => x"1800",
    100 => x"C000",
    others => x"0000"
  );

begin
  q <= rom(to_integer(unsigned(address)));
end architecture;
